library verilog;
use verilog.vl_types.all;
entity statemachine_tb is
end statemachine_tb;
