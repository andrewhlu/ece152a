library verilog;
use verilog.vl_types.all;
entity test_tb is
end test_tb;
