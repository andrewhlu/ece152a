library verilog;
use verilog.vl_types.all;
entity big_number_first_tb is
end big_number_first_tb;
