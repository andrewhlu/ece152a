library verilog;
use verilog.vl_types.all;
entity lab1_top_tb is
end lab1_top_tb;
