library verilog;
use verilog.vl_types.all;
entity float_add_tb is
end float_add_tb;
