library verilog;
use verilog.vl_types.all;
entity shifter_tb is
end shifter_tb;
