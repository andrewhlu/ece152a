library verilog;
use verilog.vl_types.all;
entity lab2_fa_tb is
end lab2_fa_tb;
