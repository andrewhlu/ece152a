library verilog;
use verilog.vl_types.all;
entity lab2_2ba_tb is
end lab2_2ba_tb;
