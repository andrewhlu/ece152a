library verilog;
use verilog.vl_types.all;
entity lab2_4ba2_tb is
end lab2_4ba2_tb;
